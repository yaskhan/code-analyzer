module parsers

import regex

pub struct KotlinParser {}

pub fn (p KotlinParser) get_extensions() []string {
	return ['.kt', '.kts']
}

pub fn (p KotlinParser) parse(content string, file_path string) ParseResult {
	mut result := ParseResult{
		file_path: file_path
		elements:  []CodeElement{}
	}

	lines := content.split_into_lines()

	for i, line in lines {
		trimmed := line.trim_space()

		// Skip empty lines
		if trimmed.len == 0 {
			continue
		}

		// Parse class definitions
		if trimmed.starts_with('class ') || trimmed.starts_with('data class ')
			|| trimmed.starts_with('object ') || trimmed.starts_with('interface ') {
			result.elements << p.parse_class(lines, i)
		}
		// Parse function/method definitions
		else if trimmed.starts_with('fun ') {
			element := p.parse_function(lines, i)
			if element.name != '' {
				result.elements << element
			}
		}
	}

	return result
}

fn (p KotlinParser) parse_class(lines []string, idx int) CodeElement {
	line := lines[idx].trim_space()

	mut class_name := ''
	mut parent := ''
	mut element_type := 'class'

	// Determine element type and extract class name
	if line.starts_with('data class ') {
		element_type = 'data class'
		mut re := regex.regex_opt(r'data\s+class\s+(\w+)') or { panic(err) }
		start, _ := re.match_string(line)
		if start >= 0 {
			groups := re.get_group_list()
			if groups.len > 0 {
				class_name = line[groups[0].start..groups[0].end]
			}
		}
	} else if line.starts_with('interface ') {
		element_type = 'interface'
		mut re := regex.regex_opt(r'interface\s+(\w+)') or { panic(err) }
		start, _ := re.match_string(line)
		if start >= 0 {
			groups := re.get_group_list()
			if groups.len > 0 {
				class_name = line[groups[0].start..groups[0].end]
			}
		}
	} else if line.starts_with('object ') {
		element_type = 'object'
		mut re := regex.regex_opt(r'object\s+(\w+)') or { panic(err) }
		start, _ := re.match_string(line)
		if start >= 0 {
			groups := re.get_group_list()
			if groups.len > 0 {
				class_name = line[groups[0].start..groups[0].end]
			}
		}
	} else {
		// Regular class
		mut re := regex.regex_opt(r'class\s+(\w+)') or { panic(err) }
		start, _ := re.match_string(line)
		if start >= 0 {
			groups := re.get_group_list()
			if groups.len > 0 {
				class_name = line[groups[0].start..groups[0].end]
			}
		}
	}

	// Extract parent class from inheritance (after colon)
	mut extends_re := regex.regex_opt(r':\s*([\w\s,]+)') or { panic(err) }
	extends_start, _ := extends_re.match_string(line)
	if extends_start >= 0 {
		extends_groups := extends_re.get_group_list()
		if extends_groups.len > 0 {
			parent = line[extends_groups[0].start..extends_groups[0].end].split(',')[0].trim_space()
		}
	}

	doc := extract_doc_lines(lines, idx, 5)

	return CodeElement{
		element_type: element_type
		name:         class_name
		parent:       parent
		doc:          doc
		line_number:  idx + 1
	}
}

fn (p KotlinParser) parse_function(lines []string, idx int) CodeElement {
	line := lines[idx].trim_space()

	mut func_name := ''
	mut access := 'public'

	// Check for access modifiers before 'fun'
	if line.starts_with('private fun ') {
		access = 'private'
	} else if line.starts_with('protected fun ') {
		access = 'protected'
	} else if line.starts_with('internal fun ') {
		access = 'internal'
	}

	// Extract function name
	mut re := regex.regex_opt(r'fun\s+(\w+)\s*\(') or { panic(err) }
	start, _ := re.match_string(line)

	if start >= 0 {
		groups := re.get_group_list()
		if groups.len > 0 {
			func_name = line[groups[0].start..groups[0].end]
		}
	}

	doc := extract_doc_lines(lines, idx, 2)

	// Determine if it's a method or function based on indentation
	element_type := if lines[idx].starts_with(' ') || lines[idx].starts_with('\t') {
		'method'
	} else {
		'function'
	}

	return CodeElement{
		element_type: element_type
		name:         func_name
		access:       access
		doc:          doc
		line_number:  idx + 1
	}
}
